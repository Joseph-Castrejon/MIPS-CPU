module and(a,b,q);
input a,b;
ouput q;


assign q = a & b;

endmodule